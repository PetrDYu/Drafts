
module nios2test (
	clk_clk,
	gpio_export,
	reset_reset_n);	

	input		clk_clk;
	output	[9:0]	gpio_export;
	input		reset_reset_n;
endmodule
