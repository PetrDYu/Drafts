// oscill_nios.v

// Generated using ACDS version 16.0 211

`timescale 1 ps / 1 ps
module oscill_nios (
		input  wire       audio_ADCDAT,                         //                         audio.ADCDAT
		input  wire       audio_ADCLRCK,                        //                              .ADCLRCK
		input  wire       audio_BCLK,                           //                              .BCLK
		output wire       audio_DACDAT,                         //                              .DACDAT
		input  wire       audio_DACLRCK,                        //                              .DACLRCK
		output wire       audio_clk_clk,                        //                     audio_clk.clk
		inout  wire       audio_config_SDAT,                    //                  audio_config.SDAT
		output wire       audio_config_SCLK,                    //                              .SCLK
		input  wire       clk_clk,                              //                           clk.clk
		output wire [6:0] pio_hex_0_external_connection_export, // pio_hex_0_external_connection.export
		output wire [6:0] pio_hex_1_external_connection_export, // pio_hex_1_external_connection.export
		output wire [6:0] pio_hex_2_external_connection_export, // pio_hex_2_external_connection.export
		output wire [6:0] pio_hex_3_external_connection_export, // pio_hex_3_external_connection.export
		output wire [6:0] pio_hex_4_external_connection_export, // pio_hex_4_external_connection.export
		output wire [6:0] pio_hex_5_external_connection_export, // pio_hex_5_external_connection.export
		input  wire [2:0] pio_key_external_connection_export,   //   pio_key_external_connection.export
		output wire [9:0] pio_led_external_connection_export,   //   pio_led_external_connection.export
		input  wire [9:0] pio_sw_external_connection_export,    //    pio_sw_external_connection.export
		input  wire       reset_reset_n,                        //                         reset.reset_n
		output wire       vga_CLK,                              //                           vga.CLK
		output wire       vga_HS,                               //                              .HS
		output wire       vga_VS,                               //                              .VS
		output wire       vga_BLANK,                            //                              .BLANK
		output wire       vga_SYNC,                             //                              .SYNC
		output wire [7:0] vga_R,                                //                              .R
		output wire [7:0] vga_G,                                //                              .G
		output wire [7:0] vga_B                                 //                              .B
	);

	wire         video_dual_clock_buffer_avalon_dc_buffer_source_valid;                      // video_dual_clock_buffer:stream_out_valid -> vga_contr:valid
	wire  [29:0] video_dual_clock_buffer_avalon_dc_buffer_source_data;                       // video_dual_clock_buffer:stream_out_data -> vga_contr:data
	wire         video_dual_clock_buffer_avalon_dc_buffer_source_ready;                      // vga_contr:ready -> video_dual_clock_buffer:stream_out_ready
	wire         video_dual_clock_buffer_avalon_dc_buffer_source_startofpacket;              // video_dual_clock_buffer:stream_out_startofpacket -> vga_contr:startofpacket
	wire         video_dual_clock_buffer_avalon_dc_buffer_source_endofpacket;                // video_dual_clock_buffer:stream_out_endofpacket -> vga_contr:endofpacket
	wire         video_pixel_buffer_dma_0_avalon_pixel_source_valid;                         // video_pixel_buffer_dma_0:stream_valid -> video_rgb_resampler_0:stream_in_valid
	wire   [7:0] video_pixel_buffer_dma_0_avalon_pixel_source_data;                          // video_pixel_buffer_dma_0:stream_data -> video_rgb_resampler_0:stream_in_data
	wire         video_pixel_buffer_dma_0_avalon_pixel_source_ready;                         // video_rgb_resampler_0:stream_in_ready -> video_pixel_buffer_dma_0:stream_ready
	wire         video_pixel_buffer_dma_0_avalon_pixel_source_startofpacket;                 // video_pixel_buffer_dma_0:stream_startofpacket -> video_rgb_resampler_0:stream_in_startofpacket
	wire         video_pixel_buffer_dma_0_avalon_pixel_source_endofpacket;                   // video_pixel_buffer_dma_0:stream_endofpacket -> video_rgb_resampler_0:stream_in_endofpacket
	wire         video_rgb_resampler_0_avalon_rgb_source_valid;                              // video_rgb_resampler_0:stream_out_valid -> video_scaler_0:stream_in_valid
	wire  [29:0] video_rgb_resampler_0_avalon_rgb_source_data;                               // video_rgb_resampler_0:stream_out_data -> video_scaler_0:stream_in_data
	wire         video_rgb_resampler_0_avalon_rgb_source_ready;                              // video_scaler_0:stream_in_ready -> video_rgb_resampler_0:stream_out_ready
	wire         video_rgb_resampler_0_avalon_rgb_source_startofpacket;                      // video_rgb_resampler_0:stream_out_startofpacket -> video_scaler_0:stream_in_startofpacket
	wire         video_rgb_resampler_0_avalon_rgb_source_endofpacket;                        // video_rgb_resampler_0:stream_out_endofpacket -> video_scaler_0:stream_in_endofpacket
	wire         video_scaler_0_avalon_scaler_source_valid;                                  // video_scaler_0:stream_out_valid -> video_dual_clock_buffer:stream_in_valid
	wire  [29:0] video_scaler_0_avalon_scaler_source_data;                                   // video_scaler_0:stream_out_data -> video_dual_clock_buffer:stream_in_data
	wire         video_scaler_0_avalon_scaler_source_ready;                                  // video_dual_clock_buffer:stream_in_ready -> video_scaler_0:stream_out_ready
	wire         video_scaler_0_avalon_scaler_source_startofpacket;                          // video_scaler_0:stream_out_startofpacket -> video_dual_clock_buffer:stream_in_startofpacket
	wire         video_scaler_0_avalon_scaler_source_endofpacket;                            // video_scaler_0:stream_out_endofpacket -> video_dual_clock_buffer:stream_in_endofpacket
	wire         pll_vga_outclk0_clk;                                                        // pll_vga:outclk_0 -> [rst_controller_002:clk, vga_contr:clk, video_dual_clock_buffer:clk_stream_out]
	wire         video_pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest;               // mm_interconnect_0:video_pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest -> video_pixel_buffer_dma_0:master_waitrequest
	wire   [7:0] video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdata;                  // mm_interconnect_0:video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdata -> video_pixel_buffer_dma_0:master_readdata
	wire  [31:0] video_pixel_buffer_dma_0_avalon_pixel_dma_master_address;                   // video_pixel_buffer_dma_0:master_address -> mm_interconnect_0:video_pixel_buffer_dma_0_avalon_pixel_dma_master_address
	wire         video_pixel_buffer_dma_0_avalon_pixel_dma_master_read;                      // video_pixel_buffer_dma_0:master_read -> mm_interconnect_0:video_pixel_buffer_dma_0_avalon_pixel_dma_master_read
	wire         video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid;             // mm_interconnect_0:video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid -> video_pixel_buffer_dma_0:master_readdatavalid
	wire         video_pixel_buffer_dma_0_avalon_pixel_dma_master_lock;                      // video_pixel_buffer_dma_0:master_arbiterlock -> mm_interconnect_0:video_pixel_buffer_dma_0_avalon_pixel_dma_master_lock
	wire  [31:0] niosii_data_master_readdata;                                                // mm_interconnect_0:niosII_data_master_readdata -> niosII:d_readdata
	wire         niosii_data_master_waitrequest;                                             // mm_interconnect_0:niosII_data_master_waitrequest -> niosII:d_waitrequest
	wire         niosii_data_master_debugaccess;                                             // niosII:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:niosII_data_master_debugaccess
	wire  [20:0] niosii_data_master_address;                                                 // niosII:d_address -> mm_interconnect_0:niosII_data_master_address
	wire   [3:0] niosii_data_master_byteenable;                                              // niosII:d_byteenable -> mm_interconnect_0:niosII_data_master_byteenable
	wire         niosii_data_master_read;                                                    // niosII:d_read -> mm_interconnect_0:niosII_data_master_read
	wire         niosii_data_master_readdatavalid;                                           // mm_interconnect_0:niosII_data_master_readdatavalid -> niosII:d_readdatavalid
	wire         niosii_data_master_write;                                                   // niosII:d_write -> mm_interconnect_0:niosII_data_master_write
	wire  [31:0] niosii_data_master_writedata;                                               // niosII:d_writedata -> mm_interconnect_0:niosII_data_master_writedata
	wire  [31:0] niosii_instruction_master_readdata;                                         // mm_interconnect_0:niosII_instruction_master_readdata -> niosII:i_readdata
	wire         niosii_instruction_master_waitrequest;                                      // mm_interconnect_0:niosII_instruction_master_waitrequest -> niosII:i_waitrequest
	wire  [20:0] niosii_instruction_master_address;                                          // niosII:i_address -> mm_interconnect_0:niosII_instruction_master_address
	wire         niosii_instruction_master_read;                                             // niosII:i_read -> mm_interconnect_0:niosII_instruction_master_read
	wire         niosii_instruction_master_readdatavalid;                                    // mm_interconnect_0:niosII_instruction_master_readdatavalid -> niosII:i_readdatavalid
	wire  [31:0] mm_interconnect_0_niosii_debug_mem_slave_readdata;                          // niosII:debug_mem_slave_readdata -> mm_interconnect_0:niosII_debug_mem_slave_readdata
	wire         mm_interconnect_0_niosii_debug_mem_slave_waitrequest;                       // niosII:debug_mem_slave_waitrequest -> mm_interconnect_0:niosII_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_niosii_debug_mem_slave_debugaccess;                       // mm_interconnect_0:niosII_debug_mem_slave_debugaccess -> niosII:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_niosii_debug_mem_slave_address;                           // mm_interconnect_0:niosII_debug_mem_slave_address -> niosII:debug_mem_slave_address
	wire         mm_interconnect_0_niosii_debug_mem_slave_read;                              // mm_interconnect_0:niosII_debug_mem_slave_read -> niosII:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_niosii_debug_mem_slave_byteenable;                        // mm_interconnect_0:niosII_debug_mem_slave_byteenable -> niosII:debug_mem_slave_byteenable
	wire         mm_interconnect_0_niosii_debug_mem_slave_write;                             // mm_interconnect_0:niosII_debug_mem_slave_write -> niosII:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_niosii_debug_mem_slave_writedata;                         // mm_interconnect_0:niosII_debug_mem_slave_writedata -> niosII:debug_mem_slave_writedata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;                   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;                     // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;                  // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;                      // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                         // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;                    // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire         mm_interconnect_0_onchip_memory_s1_chipselect;                              // mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_readdata;                                // onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	wire  [16:0] mm_interconnect_0_onchip_memory_s1_address;                                 // mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	wire   [3:0] mm_interconnect_0_onchip_memory_s1_byteenable;                              // mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	wire         mm_interconnect_0_onchip_memory_s1_write;                                   // mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_writedata;                               // mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	wire         mm_interconnect_0_onchip_memory_s1_clken;                                   // mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	wire         mm_interconnect_0_audio_transf_avalon_audio_slave_chipselect;               // mm_interconnect_0:audio_transf_avalon_audio_slave_chipselect -> audio_transf:chipselect
	wire  [31:0] mm_interconnect_0_audio_transf_avalon_audio_slave_readdata;                 // audio_transf:readdata -> mm_interconnect_0:audio_transf_avalon_audio_slave_readdata
	wire   [1:0] mm_interconnect_0_audio_transf_avalon_audio_slave_address;                  // mm_interconnect_0:audio_transf_avalon_audio_slave_address -> audio_transf:address
	wire         mm_interconnect_0_audio_transf_avalon_audio_slave_read;                     // mm_interconnect_0:audio_transf_avalon_audio_slave_read -> audio_transf:read
	wire         mm_interconnect_0_audio_transf_avalon_audio_slave_write;                    // mm_interconnect_0:audio_transf_avalon_audio_slave_write -> audio_transf:write
	wire  [31:0] mm_interconnect_0_audio_transf_avalon_audio_slave_writedata;                // mm_interconnect_0:audio_transf_avalon_audio_slave_writedata -> audio_transf:writedata
	wire  [31:0] mm_interconnect_0_av_config_avalon_av_config_slave_readdata;                // av_config:readdata -> mm_interconnect_0:av_config_avalon_av_config_slave_readdata
	wire         mm_interconnect_0_av_config_avalon_av_config_slave_waitrequest;             // av_config:waitrequest -> mm_interconnect_0:av_config_avalon_av_config_slave_waitrequest
	wire   [1:0] mm_interconnect_0_av_config_avalon_av_config_slave_address;                 // mm_interconnect_0:av_config_avalon_av_config_slave_address -> av_config:address
	wire         mm_interconnect_0_av_config_avalon_av_config_slave_read;                    // mm_interconnect_0:av_config_avalon_av_config_slave_read -> av_config:read
	wire   [3:0] mm_interconnect_0_av_config_avalon_av_config_slave_byteenable;              // mm_interconnect_0:av_config_avalon_av_config_slave_byteenable -> av_config:byteenable
	wire         mm_interconnect_0_av_config_avalon_av_config_slave_write;                   // mm_interconnect_0:av_config_avalon_av_config_slave_write -> av_config:write
	wire  [31:0] mm_interconnect_0_av_config_avalon_av_config_slave_writedata;               // mm_interconnect_0:av_config_avalon_av_config_slave_writedata -> av_config:writedata
	wire  [31:0] mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_readdata;   // video_pixel_buffer_dma_0:slave_readdata -> mm_interconnect_0:video_pixel_buffer_dma_0_avalon_control_slave_readdata
	wire   [1:0] mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_address;    // mm_interconnect_0:video_pixel_buffer_dma_0_avalon_control_slave_address -> video_pixel_buffer_dma_0:slave_address
	wire         mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_read;       // mm_interconnect_0:video_pixel_buffer_dma_0_avalon_control_slave_read -> video_pixel_buffer_dma_0:slave_read
	wire   [3:0] mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_byteenable; // mm_interconnect_0:video_pixel_buffer_dma_0_avalon_control_slave_byteenable -> video_pixel_buffer_dma_0:slave_byteenable
	wire         mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_write;      // mm_interconnect_0:video_pixel_buffer_dma_0_avalon_control_slave_write -> video_pixel_buffer_dma_0:slave_write
	wire  [31:0] mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_writedata;  // mm_interconnect_0:video_pixel_buffer_dma_0_avalon_control_slave_writedata -> video_pixel_buffer_dma_0:slave_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_control_slave_readdata;                        // sysid_qsys:readdata -> mm_interconnect_0:sysid_qsys_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_control_slave_address;                         // mm_interconnect_0:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire  [31:0] mm_interconnect_0_pio_key_s1_readdata;                                      // pio_key:readdata -> mm_interconnect_0:pio_key_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_key_s1_address;                                       // mm_interconnect_0:pio_key_s1_address -> pio_key:address
	wire         mm_interconnect_0_pio_led_s1_chipselect;                                    // mm_interconnect_0:pio_led_s1_chipselect -> pio_led:chipselect
	wire  [31:0] mm_interconnect_0_pio_led_s1_readdata;                                      // pio_led:readdata -> mm_interconnect_0:pio_led_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_led_s1_address;                                       // mm_interconnect_0:pio_led_s1_address -> pio_led:address
	wire         mm_interconnect_0_pio_led_s1_write;                                         // mm_interconnect_0:pio_led_s1_write -> pio_led:write_n
	wire  [31:0] mm_interconnect_0_pio_led_s1_writedata;                                     // mm_interconnect_0:pio_led_s1_writedata -> pio_led:writedata
	wire         mm_interconnect_0_pio_hex_0_s1_chipselect;                                  // mm_interconnect_0:pio_hex_0_s1_chipselect -> pio_hex_0:chipselect
	wire  [31:0] mm_interconnect_0_pio_hex_0_s1_readdata;                                    // pio_hex_0:readdata -> mm_interconnect_0:pio_hex_0_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_hex_0_s1_address;                                     // mm_interconnect_0:pio_hex_0_s1_address -> pio_hex_0:address
	wire         mm_interconnect_0_pio_hex_0_s1_write;                                       // mm_interconnect_0:pio_hex_0_s1_write -> pio_hex_0:write_n
	wire  [31:0] mm_interconnect_0_pio_hex_0_s1_writedata;                                   // mm_interconnect_0:pio_hex_0_s1_writedata -> pio_hex_0:writedata
	wire  [31:0] mm_interconnect_0_pio_sw_s1_readdata;                                       // pio_sw:readdata -> mm_interconnect_0:pio_sw_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_sw_s1_address;                                        // mm_interconnect_0:pio_sw_s1_address -> pio_sw:address
	wire         mm_interconnect_0_pio_hex_1_s1_chipselect;                                  // mm_interconnect_0:pio_hex_1_s1_chipselect -> pio_hex_1:chipselect
	wire  [31:0] mm_interconnect_0_pio_hex_1_s1_readdata;                                    // pio_hex_1:readdata -> mm_interconnect_0:pio_hex_1_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_hex_1_s1_address;                                     // mm_interconnect_0:pio_hex_1_s1_address -> pio_hex_1:address
	wire         mm_interconnect_0_pio_hex_1_s1_write;                                       // mm_interconnect_0:pio_hex_1_s1_write -> pio_hex_1:write_n
	wire  [31:0] mm_interconnect_0_pio_hex_1_s1_writedata;                                   // mm_interconnect_0:pio_hex_1_s1_writedata -> pio_hex_1:writedata
	wire         mm_interconnect_0_pio_hex_2_s1_chipselect;                                  // mm_interconnect_0:pio_hex_2_s1_chipselect -> pio_hex_2:chipselect
	wire  [31:0] mm_interconnect_0_pio_hex_2_s1_readdata;                                    // pio_hex_2:readdata -> mm_interconnect_0:pio_hex_2_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_hex_2_s1_address;                                     // mm_interconnect_0:pio_hex_2_s1_address -> pio_hex_2:address
	wire         mm_interconnect_0_pio_hex_2_s1_write;                                       // mm_interconnect_0:pio_hex_2_s1_write -> pio_hex_2:write_n
	wire  [31:0] mm_interconnect_0_pio_hex_2_s1_writedata;                                   // mm_interconnect_0:pio_hex_2_s1_writedata -> pio_hex_2:writedata
	wire         mm_interconnect_0_pio_hex_3_s1_chipselect;                                  // mm_interconnect_0:pio_hex_3_s1_chipselect -> pio_hex_3:chipselect
	wire  [31:0] mm_interconnect_0_pio_hex_3_s1_readdata;                                    // pio_hex_3:readdata -> mm_interconnect_0:pio_hex_3_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_hex_3_s1_address;                                     // mm_interconnect_0:pio_hex_3_s1_address -> pio_hex_3:address
	wire         mm_interconnect_0_pio_hex_3_s1_write;                                       // mm_interconnect_0:pio_hex_3_s1_write -> pio_hex_3:write_n
	wire  [31:0] mm_interconnect_0_pio_hex_3_s1_writedata;                                   // mm_interconnect_0:pio_hex_3_s1_writedata -> pio_hex_3:writedata
	wire         mm_interconnect_0_pio_hex_4_s1_chipselect;                                  // mm_interconnect_0:pio_hex_4_s1_chipselect -> pio_hex_4:chipselect
	wire  [31:0] mm_interconnect_0_pio_hex_4_s1_readdata;                                    // pio_hex_4:readdata -> mm_interconnect_0:pio_hex_4_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_hex_4_s1_address;                                     // mm_interconnect_0:pio_hex_4_s1_address -> pio_hex_4:address
	wire         mm_interconnect_0_pio_hex_4_s1_write;                                       // mm_interconnect_0:pio_hex_4_s1_write -> pio_hex_4:write_n
	wire  [31:0] mm_interconnect_0_pio_hex_4_s1_writedata;                                   // mm_interconnect_0:pio_hex_4_s1_writedata -> pio_hex_4:writedata
	wire         mm_interconnect_0_pio_hex_5_s1_chipselect;                                  // mm_interconnect_0:pio_hex_5_s1_chipselect -> pio_hex_5:chipselect
	wire  [31:0] mm_interconnect_0_pio_hex_5_s1_readdata;                                    // pio_hex_5:readdata -> mm_interconnect_0:pio_hex_5_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_hex_5_s1_address;                                     // mm_interconnect_0:pio_hex_5_s1_address -> pio_hex_5:address
	wire         mm_interconnect_0_pio_hex_5_s1_write;                                       // mm_interconnect_0:pio_hex_5_s1_write -> pio_hex_5:write_n
	wire  [31:0] mm_interconnect_0_pio_hex_5_s1_writedata;                                   // mm_interconnect_0:pio_hex_5_s1_writedata -> pio_hex_5:writedata
	wire         irq_mapper_receiver0_irq;                                                   // audio_transf:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                   // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire  [31:0] niosii_irq_irq;                                                             // irq_mapper:sender_irq -> niosII:irq
	wire         rst_controller_reset_out_reset;                                             // rst_controller:reset_out -> [audio_transf:reset, mm_interconnect_0:audio_transf_reset_reset_bridge_in_reset_reset]
	wire         audio_pll_reset_source_reset;                                               // audio_pll:reset_source_reset -> rst_controller:reset_in0
	wire         rst_controller_001_reset_out_reset;                                         // rst_controller_001:reset_out -> [av_config:reset, irq_mapper:reset, jtag_uart:rst_n, mm_interconnect_0:video_pixel_buffer_dma_0_reset_reset_bridge_in_reset_reset, niosII:reset_n, onchip_memory:reset, pio_hex_0:reset_n, pio_hex_1:reset_n, pio_hex_2:reset_n, pio_hex_3:reset_n, pio_hex_4:reset_n, pio_hex_5:reset_n, pio_key:reset_n, pio_led:reset_n, pio_sw:reset_n, rst_translator:in_reset, sysid_qsys:reset_n, video_dual_clock_buffer:reset_stream_in, video_pixel_buffer_dma_0:reset, video_rgb_resampler_0:reset, video_scaler_0:reset]
	wire         rst_controller_001_reset_out_reset_req;                                     // rst_controller_001:reset_req -> [niosII:reset_req, onchip_memory:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_002_reset_out_reset;                                         // rst_controller_002:reset_out -> [vga_contr:reset, video_dual_clock_buffer:reset_stream_out]

	oscill_nios_audio_pll audio_pll (
		.ref_clk_clk        (clk_clk),                      //      ref_clk.clk
		.ref_reset_reset    (~reset_reset_n),               //    ref_reset.reset
		.audio_clk_clk      (audio_clk_clk),                //    audio_clk.clk
		.reset_source_reset (audio_pll_reset_source_reset)  // reset_source.reset
	);

	oscill_nios_audio_transf audio_transf (
		.clk         (clk_clk),                                                      //                clk.clk
		.reset       (rst_controller_reset_out_reset),                               //              reset.reset
		.address     (mm_interconnect_0_audio_transf_avalon_audio_slave_address),    // avalon_audio_slave.address
		.chipselect  (mm_interconnect_0_audio_transf_avalon_audio_slave_chipselect), //                   .chipselect
		.read        (mm_interconnect_0_audio_transf_avalon_audio_slave_read),       //                   .read
		.write       (mm_interconnect_0_audio_transf_avalon_audio_slave_write),      //                   .write
		.writedata   (mm_interconnect_0_audio_transf_avalon_audio_slave_writedata),  //                   .writedata
		.readdata    (mm_interconnect_0_audio_transf_avalon_audio_slave_readdata),   //                   .readdata
		.irq         (irq_mapper_receiver0_irq),                                     //          interrupt.irq
		.AUD_ADCDAT  (audio_ADCDAT),                                                 // external_interface.export
		.AUD_ADCLRCK (audio_ADCLRCK),                                                //                   .export
		.AUD_BCLK    (audio_BCLK),                                                   //                   .export
		.AUD_DACDAT  (audio_DACDAT),                                                 //                   .export
		.AUD_DACLRCK (audio_DACLRCK)                                                 //                   .export
	);

	oscill_nios_av_config av_config (
		.clk         (clk_clk),                                                        //                    clk.clk
		.reset       (rst_controller_001_reset_out_reset),                             //                  reset.reset
		.address     (mm_interconnect_0_av_config_avalon_av_config_slave_address),     // avalon_av_config_slave.address
		.byteenable  (mm_interconnect_0_av_config_avalon_av_config_slave_byteenable),  //                       .byteenable
		.read        (mm_interconnect_0_av_config_avalon_av_config_slave_read),        //                       .read
		.write       (mm_interconnect_0_av_config_avalon_av_config_slave_write),       //                       .write
		.writedata   (mm_interconnect_0_av_config_avalon_av_config_slave_writedata),   //                       .writedata
		.readdata    (mm_interconnect_0_av_config_avalon_av_config_slave_readdata),    //                       .readdata
		.waitrequest (mm_interconnect_0_av_config_avalon_av_config_slave_waitrequest), //                       .waitrequest
		.I2C_SDAT    (audio_config_SDAT),                                              //     external_interface.export
		.I2C_SCLK    (audio_config_SCLK)                                               //                       .export
	);

	oscill_nios_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
	);

	oscill_nios_niosII niosii (
		.clk                                 (clk_clk),                                              //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                  //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),               //                          .reset_req
		.d_address                           (niosii_data_master_address),                           //               data_master.address
		.d_byteenable                        (niosii_data_master_byteenable),                        //                          .byteenable
		.d_read                              (niosii_data_master_read),                              //                          .read
		.d_readdata                          (niosii_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (niosii_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (niosii_data_master_write),                             //                          .write
		.d_writedata                         (niosii_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (niosii_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (niosii_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (niosii_instruction_master_address),                    //        instruction_master.address
		.i_read                              (niosii_instruction_master_read),                       //                          .read
		.i_readdata                          (niosii_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (niosii_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (niosii_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (niosii_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_niosii_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_niosii_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_niosii_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_niosii_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_niosii_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_niosii_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_niosii_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_niosii_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                      // custom_instruction_master.readra
	);

	oscill_nios_onchip_memory onchip_memory (
		.clk        (clk_clk),                                       //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),            // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req)         //       .reset_req
	);

	oscill_nios_pio_hex_0 pio_hex_0 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_pio_hex_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_hex_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_hex_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_hex_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_hex_0_s1_readdata),   //                    .readdata
		.out_port   (pio_hex_0_external_connection_export)       // external_connection.export
	);

	oscill_nios_pio_hex_0 pio_hex_1 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_pio_hex_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_hex_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_hex_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_hex_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_hex_1_s1_readdata),   //                    .readdata
		.out_port   (pio_hex_1_external_connection_export)       // external_connection.export
	);

	oscill_nios_pio_hex_0 pio_hex_2 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_pio_hex_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_hex_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_hex_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_hex_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_hex_2_s1_readdata),   //                    .readdata
		.out_port   (pio_hex_2_external_connection_export)       // external_connection.export
	);

	oscill_nios_pio_hex_0 pio_hex_3 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_pio_hex_3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_hex_3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_hex_3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_hex_3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_hex_3_s1_readdata),   //                    .readdata
		.out_port   (pio_hex_3_external_connection_export)       // external_connection.export
	);

	oscill_nios_pio_hex_0 pio_hex_4 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_pio_hex_4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_hex_4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_hex_4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_hex_4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_hex_4_s1_readdata),   //                    .readdata
		.out_port   (pio_hex_4_external_connection_export)       // external_connection.export
	);

	oscill_nios_pio_hex_0 pio_hex_5 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_pio_hex_5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_hex_5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_hex_5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_hex_5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_hex_5_s1_readdata),   //                    .readdata
		.out_port   (pio_hex_5_external_connection_export)       // external_connection.export
	);

	oscill_nios_pio_key pio_key (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),   //               reset.reset_n
		.address  (mm_interconnect_0_pio_key_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_key_s1_readdata), //                    .readdata
		.in_port  (pio_key_external_connection_export)     // external_connection.export
	);

	oscill_nios_pio_led pio_led (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_pio_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_led_s1_readdata),   //                    .readdata
		.out_port   (pio_led_external_connection_export)       // external_connection.export
	);

	oscill_nios_pio_sw pio_sw (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),  //               reset.reset_n
		.address  (mm_interconnect_0_pio_sw_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_sw_s1_readdata), //                    .readdata
		.in_port  (pio_sw_external_connection_export)     // external_connection.export
	);

	oscill_nios_pll_vga pll_vga (
		.refclk   (clk_clk),             //  refclk.clk
		.rst      (~reset_reset_n),      //   reset.reset
		.outclk_0 (pll_vga_outclk0_clk), // outclk0.clk
		.locked   ()                     // (terminated)
	);

	oscill_nios_sysid_qsys sysid_qsys (
		.clock    (clk_clk),                                             //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                 //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_control_slave_address)   //              .address
	);

	oscill_nios_vga_contr vga_contr (
		.clk           (pll_vga_outclk0_clk),                                           //                clk.clk
		.reset         (rst_controller_002_reset_out_reset),                            //              reset.reset
		.data          (video_dual_clock_buffer_avalon_dc_buffer_source_data),          //    avalon_vga_sink.data
		.startofpacket (video_dual_clock_buffer_avalon_dc_buffer_source_startofpacket), //                   .startofpacket
		.endofpacket   (video_dual_clock_buffer_avalon_dc_buffer_source_endofpacket),   //                   .endofpacket
		.valid         (video_dual_clock_buffer_avalon_dc_buffer_source_valid),         //                   .valid
		.ready         (video_dual_clock_buffer_avalon_dc_buffer_source_ready),         //                   .ready
		.VGA_CLK       (vga_CLK),                                                       // external_interface.export
		.VGA_HS        (vga_HS),                                                        //                   .export
		.VGA_VS        (vga_VS),                                                        //                   .export
		.VGA_BLANK     (vga_BLANK),                                                     //                   .export
		.VGA_SYNC      (vga_SYNC),                                                      //                   .export
		.VGA_R         (vga_R),                                                         //                   .export
		.VGA_G         (vga_G),                                                         //                   .export
		.VGA_B         (vga_B)                                                          //                   .export
	);

	oscill_nios_video_dual_clock_buffer video_dual_clock_buffer (
		.clk_stream_in            (clk_clk),                                                       //         clock_stream_in.clk
		.reset_stream_in          (rst_controller_001_reset_out_reset),                            //         reset_stream_in.reset
		.clk_stream_out           (pll_vga_outclk0_clk),                                           //        clock_stream_out.clk
		.reset_stream_out         (rst_controller_002_reset_out_reset),                            //        reset_stream_out.reset
		.stream_in_ready          (video_scaler_0_avalon_scaler_source_ready),                     //   avalon_dc_buffer_sink.ready
		.stream_in_startofpacket  (video_scaler_0_avalon_scaler_source_startofpacket),             //                        .startofpacket
		.stream_in_endofpacket    (video_scaler_0_avalon_scaler_source_endofpacket),               //                        .endofpacket
		.stream_in_valid          (video_scaler_0_avalon_scaler_source_valid),                     //                        .valid
		.stream_in_data           (video_scaler_0_avalon_scaler_source_data),                      //                        .data
		.stream_out_ready         (video_dual_clock_buffer_avalon_dc_buffer_source_ready),         // avalon_dc_buffer_source.ready
		.stream_out_startofpacket (video_dual_clock_buffer_avalon_dc_buffer_source_startofpacket), //                        .startofpacket
		.stream_out_endofpacket   (video_dual_clock_buffer_avalon_dc_buffer_source_endofpacket),   //                        .endofpacket
		.stream_out_valid         (video_dual_clock_buffer_avalon_dc_buffer_source_valid),         //                        .valid
		.stream_out_data          (video_dual_clock_buffer_avalon_dc_buffer_source_data)           //                        .data
	);

	oscill_nios_video_pixel_buffer_dma_0 video_pixel_buffer_dma_0 (
		.clk                  (clk_clk),                                                                    //                     clk.clk
		.reset                (rst_controller_001_reset_out_reset),                                         //                   reset.reset
		.master_readdatavalid (video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid),             // avalon_pixel_dma_master.readdatavalid
		.master_waitrequest   (video_pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest),               //                        .waitrequest
		.master_address       (video_pixel_buffer_dma_0_avalon_pixel_dma_master_address),                   //                        .address
		.master_arbiterlock   (video_pixel_buffer_dma_0_avalon_pixel_dma_master_lock),                      //                        .lock
		.master_read          (video_pixel_buffer_dma_0_avalon_pixel_dma_master_read),                      //                        .read
		.master_readdata      (video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdata),                  //                        .readdata
		.slave_address        (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_address),    //    avalon_control_slave.address
		.slave_byteenable     (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_byteenable), //                        .byteenable
		.slave_read           (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_read),       //                        .read
		.slave_write          (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_write),      //                        .write
		.slave_writedata      (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_writedata),  //                        .writedata
		.slave_readdata       (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_readdata),   //                        .readdata
		.stream_ready         (video_pixel_buffer_dma_0_avalon_pixel_source_ready),                         //     avalon_pixel_source.ready
		.stream_startofpacket (video_pixel_buffer_dma_0_avalon_pixel_source_startofpacket),                 //                        .startofpacket
		.stream_endofpacket   (video_pixel_buffer_dma_0_avalon_pixel_source_endofpacket),                   //                        .endofpacket
		.stream_valid         (video_pixel_buffer_dma_0_avalon_pixel_source_valid),                         //                        .valid
		.stream_data          (video_pixel_buffer_dma_0_avalon_pixel_source_data)                           //                        .data
	);

	oscill_nios_video_rgb_resampler_0 video_rgb_resampler_0 (
		.clk                      (clk_clk),                                                    //               clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                         //             reset.reset
		.stream_in_startofpacket  (video_pixel_buffer_dma_0_avalon_pixel_source_startofpacket), //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (video_pixel_buffer_dma_0_avalon_pixel_source_endofpacket),   //                  .endofpacket
		.stream_in_valid          (video_pixel_buffer_dma_0_avalon_pixel_source_valid),         //                  .valid
		.stream_in_ready          (video_pixel_buffer_dma_0_avalon_pixel_source_ready),         //                  .ready
		.stream_in_data           (video_pixel_buffer_dma_0_avalon_pixel_source_data),          //                  .data
		.stream_out_ready         (video_rgb_resampler_0_avalon_rgb_source_ready),              // avalon_rgb_source.ready
		.stream_out_startofpacket (video_rgb_resampler_0_avalon_rgb_source_startofpacket),      //                  .startofpacket
		.stream_out_endofpacket   (video_rgb_resampler_0_avalon_rgb_source_endofpacket),        //                  .endofpacket
		.stream_out_valid         (video_rgb_resampler_0_avalon_rgb_source_valid),              //                  .valid
		.stream_out_data          (video_rgb_resampler_0_avalon_rgb_source_data)                //                  .data
	);

	oscill_nios_video_scaler_0 video_scaler_0 (
		.clk                      (clk_clk),                                               //                  clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                    //                reset.reset
		.stream_in_startofpacket  (video_rgb_resampler_0_avalon_rgb_source_startofpacket), //   avalon_scaler_sink.startofpacket
		.stream_in_endofpacket    (video_rgb_resampler_0_avalon_rgb_source_endofpacket),   //                     .endofpacket
		.stream_in_valid          (video_rgb_resampler_0_avalon_rgb_source_valid),         //                     .valid
		.stream_in_ready          (video_rgb_resampler_0_avalon_rgb_source_ready),         //                     .ready
		.stream_in_data           (video_rgb_resampler_0_avalon_rgb_source_data),          //                     .data
		.stream_out_ready         (video_scaler_0_avalon_scaler_source_ready),             // avalon_scaler_source.ready
		.stream_out_startofpacket (video_scaler_0_avalon_scaler_source_startofpacket),     //                     .startofpacket
		.stream_out_endofpacket   (video_scaler_0_avalon_scaler_source_endofpacket),       //                     .endofpacket
		.stream_out_valid         (video_scaler_0_avalon_scaler_source_valid),             //                     .valid
		.stream_out_data          (video_scaler_0_avalon_scaler_source_data)               //                     .data
	);

	oscill_nios_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                                                    (clk_clk),                                                                    //                                              clk_clk.clk
		.audio_transf_reset_reset_bridge_in_reset_reset                 (rst_controller_reset_out_reset),                                             //             audio_transf_reset_reset_bridge_in_reset.reset
		.video_pixel_buffer_dma_0_reset_reset_bridge_in_reset_reset     (rst_controller_001_reset_out_reset),                                         // video_pixel_buffer_dma_0_reset_reset_bridge_in_reset.reset
		.niosII_data_master_address                                     (niosii_data_master_address),                                                 //                                   niosII_data_master.address
		.niosII_data_master_waitrequest                                 (niosii_data_master_waitrequest),                                             //                                                     .waitrequest
		.niosII_data_master_byteenable                                  (niosii_data_master_byteenable),                                              //                                                     .byteenable
		.niosII_data_master_read                                        (niosii_data_master_read),                                                    //                                                     .read
		.niosII_data_master_readdata                                    (niosii_data_master_readdata),                                                //                                                     .readdata
		.niosII_data_master_readdatavalid                               (niosii_data_master_readdatavalid),                                           //                                                     .readdatavalid
		.niosII_data_master_write                                       (niosii_data_master_write),                                                   //                                                     .write
		.niosII_data_master_writedata                                   (niosii_data_master_writedata),                                               //                                                     .writedata
		.niosII_data_master_debugaccess                                 (niosii_data_master_debugaccess),                                             //                                                     .debugaccess
		.niosII_instruction_master_address                              (niosii_instruction_master_address),                                          //                            niosII_instruction_master.address
		.niosII_instruction_master_waitrequest                          (niosii_instruction_master_waitrequest),                                      //                                                     .waitrequest
		.niosII_instruction_master_read                                 (niosii_instruction_master_read),                                             //                                                     .read
		.niosII_instruction_master_readdata                             (niosii_instruction_master_readdata),                                         //                                                     .readdata
		.niosII_instruction_master_readdatavalid                        (niosii_instruction_master_readdatavalid),                                    //                                                     .readdatavalid
		.video_pixel_buffer_dma_0_avalon_pixel_dma_master_address       (video_pixel_buffer_dma_0_avalon_pixel_dma_master_address),                   //     video_pixel_buffer_dma_0_avalon_pixel_dma_master.address
		.video_pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest   (video_pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest),               //                                                     .waitrequest
		.video_pixel_buffer_dma_0_avalon_pixel_dma_master_read          (video_pixel_buffer_dma_0_avalon_pixel_dma_master_read),                      //                                                     .read
		.video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdata      (video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdata),                  //                                                     .readdata
		.video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid (video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid),             //                                                     .readdatavalid
		.video_pixel_buffer_dma_0_avalon_pixel_dma_master_lock          (video_pixel_buffer_dma_0_avalon_pixel_dma_master_lock),                      //                                                     .lock
		.audio_transf_avalon_audio_slave_address                        (mm_interconnect_0_audio_transf_avalon_audio_slave_address),                  //                      audio_transf_avalon_audio_slave.address
		.audio_transf_avalon_audio_slave_write                          (mm_interconnect_0_audio_transf_avalon_audio_slave_write),                    //                                                     .write
		.audio_transf_avalon_audio_slave_read                           (mm_interconnect_0_audio_transf_avalon_audio_slave_read),                     //                                                     .read
		.audio_transf_avalon_audio_slave_readdata                       (mm_interconnect_0_audio_transf_avalon_audio_slave_readdata),                 //                                                     .readdata
		.audio_transf_avalon_audio_slave_writedata                      (mm_interconnect_0_audio_transf_avalon_audio_slave_writedata),                //                                                     .writedata
		.audio_transf_avalon_audio_slave_chipselect                     (mm_interconnect_0_audio_transf_avalon_audio_slave_chipselect),               //                                                     .chipselect
		.av_config_avalon_av_config_slave_address                       (mm_interconnect_0_av_config_avalon_av_config_slave_address),                 //                     av_config_avalon_av_config_slave.address
		.av_config_avalon_av_config_slave_write                         (mm_interconnect_0_av_config_avalon_av_config_slave_write),                   //                                                     .write
		.av_config_avalon_av_config_slave_read                          (mm_interconnect_0_av_config_avalon_av_config_slave_read),                    //                                                     .read
		.av_config_avalon_av_config_slave_readdata                      (mm_interconnect_0_av_config_avalon_av_config_slave_readdata),                //                                                     .readdata
		.av_config_avalon_av_config_slave_writedata                     (mm_interconnect_0_av_config_avalon_av_config_slave_writedata),               //                                                     .writedata
		.av_config_avalon_av_config_slave_byteenable                    (mm_interconnect_0_av_config_avalon_av_config_slave_byteenable),              //                                                     .byteenable
		.av_config_avalon_av_config_slave_waitrequest                   (mm_interconnect_0_av_config_avalon_av_config_slave_waitrequest),             //                                                     .waitrequest
		.jtag_uart_avalon_jtag_slave_address                            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),                      //                          jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),                        //                                                     .write
		.jtag_uart_avalon_jtag_slave_read                               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),                         //                                                     .read
		.jtag_uart_avalon_jtag_slave_readdata                           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),                     //                                                     .readdata
		.jtag_uart_avalon_jtag_slave_writedata                          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),                    //                                                     .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),                  //                                                     .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),                   //                                                     .chipselect
		.niosII_debug_mem_slave_address                                 (mm_interconnect_0_niosii_debug_mem_slave_address),                           //                               niosII_debug_mem_slave.address
		.niosII_debug_mem_slave_write                                   (mm_interconnect_0_niosii_debug_mem_slave_write),                             //                                                     .write
		.niosII_debug_mem_slave_read                                    (mm_interconnect_0_niosii_debug_mem_slave_read),                              //                                                     .read
		.niosII_debug_mem_slave_readdata                                (mm_interconnect_0_niosii_debug_mem_slave_readdata),                          //                                                     .readdata
		.niosII_debug_mem_slave_writedata                               (mm_interconnect_0_niosii_debug_mem_slave_writedata),                         //                                                     .writedata
		.niosII_debug_mem_slave_byteenable                              (mm_interconnect_0_niosii_debug_mem_slave_byteenable),                        //                                                     .byteenable
		.niosII_debug_mem_slave_waitrequest                             (mm_interconnect_0_niosii_debug_mem_slave_waitrequest),                       //                                                     .waitrequest
		.niosII_debug_mem_slave_debugaccess                             (mm_interconnect_0_niosii_debug_mem_slave_debugaccess),                       //                                                     .debugaccess
		.onchip_memory_s1_address                                       (mm_interconnect_0_onchip_memory_s1_address),                                 //                                     onchip_memory_s1.address
		.onchip_memory_s1_write                                         (mm_interconnect_0_onchip_memory_s1_write),                                   //                                                     .write
		.onchip_memory_s1_readdata                                      (mm_interconnect_0_onchip_memory_s1_readdata),                                //                                                     .readdata
		.onchip_memory_s1_writedata                                     (mm_interconnect_0_onchip_memory_s1_writedata),                               //                                                     .writedata
		.onchip_memory_s1_byteenable                                    (mm_interconnect_0_onchip_memory_s1_byteenable),                              //                                                     .byteenable
		.onchip_memory_s1_chipselect                                    (mm_interconnect_0_onchip_memory_s1_chipselect),                              //                                                     .chipselect
		.onchip_memory_s1_clken                                         (mm_interconnect_0_onchip_memory_s1_clken),                                   //                                                     .clken
		.pio_hex_0_s1_address                                           (mm_interconnect_0_pio_hex_0_s1_address),                                     //                                         pio_hex_0_s1.address
		.pio_hex_0_s1_write                                             (mm_interconnect_0_pio_hex_0_s1_write),                                       //                                                     .write
		.pio_hex_0_s1_readdata                                          (mm_interconnect_0_pio_hex_0_s1_readdata),                                    //                                                     .readdata
		.pio_hex_0_s1_writedata                                         (mm_interconnect_0_pio_hex_0_s1_writedata),                                   //                                                     .writedata
		.pio_hex_0_s1_chipselect                                        (mm_interconnect_0_pio_hex_0_s1_chipselect),                                  //                                                     .chipselect
		.pio_hex_1_s1_address                                           (mm_interconnect_0_pio_hex_1_s1_address),                                     //                                         pio_hex_1_s1.address
		.pio_hex_1_s1_write                                             (mm_interconnect_0_pio_hex_1_s1_write),                                       //                                                     .write
		.pio_hex_1_s1_readdata                                          (mm_interconnect_0_pio_hex_1_s1_readdata),                                    //                                                     .readdata
		.pio_hex_1_s1_writedata                                         (mm_interconnect_0_pio_hex_1_s1_writedata),                                   //                                                     .writedata
		.pio_hex_1_s1_chipselect                                        (mm_interconnect_0_pio_hex_1_s1_chipselect),                                  //                                                     .chipselect
		.pio_hex_2_s1_address                                           (mm_interconnect_0_pio_hex_2_s1_address),                                     //                                         pio_hex_2_s1.address
		.pio_hex_2_s1_write                                             (mm_interconnect_0_pio_hex_2_s1_write),                                       //                                                     .write
		.pio_hex_2_s1_readdata                                          (mm_interconnect_0_pio_hex_2_s1_readdata),                                    //                                                     .readdata
		.pio_hex_2_s1_writedata                                         (mm_interconnect_0_pio_hex_2_s1_writedata),                                   //                                                     .writedata
		.pio_hex_2_s1_chipselect                                        (mm_interconnect_0_pio_hex_2_s1_chipselect),                                  //                                                     .chipselect
		.pio_hex_3_s1_address                                           (mm_interconnect_0_pio_hex_3_s1_address),                                     //                                         pio_hex_3_s1.address
		.pio_hex_3_s1_write                                             (mm_interconnect_0_pio_hex_3_s1_write),                                       //                                                     .write
		.pio_hex_3_s1_readdata                                          (mm_interconnect_0_pio_hex_3_s1_readdata),                                    //                                                     .readdata
		.pio_hex_3_s1_writedata                                         (mm_interconnect_0_pio_hex_3_s1_writedata),                                   //                                                     .writedata
		.pio_hex_3_s1_chipselect                                        (mm_interconnect_0_pio_hex_3_s1_chipselect),                                  //                                                     .chipselect
		.pio_hex_4_s1_address                                           (mm_interconnect_0_pio_hex_4_s1_address),                                     //                                         pio_hex_4_s1.address
		.pio_hex_4_s1_write                                             (mm_interconnect_0_pio_hex_4_s1_write),                                       //                                                     .write
		.pio_hex_4_s1_readdata                                          (mm_interconnect_0_pio_hex_4_s1_readdata),                                    //                                                     .readdata
		.pio_hex_4_s1_writedata                                         (mm_interconnect_0_pio_hex_4_s1_writedata),                                   //                                                     .writedata
		.pio_hex_4_s1_chipselect                                        (mm_interconnect_0_pio_hex_4_s1_chipselect),                                  //                                                     .chipselect
		.pio_hex_5_s1_address                                           (mm_interconnect_0_pio_hex_5_s1_address),                                     //                                         pio_hex_5_s1.address
		.pio_hex_5_s1_write                                             (mm_interconnect_0_pio_hex_5_s1_write),                                       //                                                     .write
		.pio_hex_5_s1_readdata                                          (mm_interconnect_0_pio_hex_5_s1_readdata),                                    //                                                     .readdata
		.pio_hex_5_s1_writedata                                         (mm_interconnect_0_pio_hex_5_s1_writedata),                                   //                                                     .writedata
		.pio_hex_5_s1_chipselect                                        (mm_interconnect_0_pio_hex_5_s1_chipselect),                                  //                                                     .chipselect
		.pio_key_s1_address                                             (mm_interconnect_0_pio_key_s1_address),                                       //                                           pio_key_s1.address
		.pio_key_s1_readdata                                            (mm_interconnect_0_pio_key_s1_readdata),                                      //                                                     .readdata
		.pio_led_s1_address                                             (mm_interconnect_0_pio_led_s1_address),                                       //                                           pio_led_s1.address
		.pio_led_s1_write                                               (mm_interconnect_0_pio_led_s1_write),                                         //                                                     .write
		.pio_led_s1_readdata                                            (mm_interconnect_0_pio_led_s1_readdata),                                      //                                                     .readdata
		.pio_led_s1_writedata                                           (mm_interconnect_0_pio_led_s1_writedata),                                     //                                                     .writedata
		.pio_led_s1_chipselect                                          (mm_interconnect_0_pio_led_s1_chipselect),                                    //                                                     .chipselect
		.pio_sw_s1_address                                              (mm_interconnect_0_pio_sw_s1_address),                                        //                                            pio_sw_s1.address
		.pio_sw_s1_readdata                                             (mm_interconnect_0_pio_sw_s1_readdata),                                       //                                                     .readdata
		.sysid_qsys_control_slave_address                               (mm_interconnect_0_sysid_qsys_control_slave_address),                         //                             sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata                              (mm_interconnect_0_sysid_qsys_control_slave_readdata),                        //                                                     .readdata
		.video_pixel_buffer_dma_0_avalon_control_slave_address          (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_address),    //        video_pixel_buffer_dma_0_avalon_control_slave.address
		.video_pixel_buffer_dma_0_avalon_control_slave_write            (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_write),      //                                                     .write
		.video_pixel_buffer_dma_0_avalon_control_slave_read             (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_read),       //                                                     .read
		.video_pixel_buffer_dma_0_avalon_control_slave_readdata         (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_readdata),   //                                                     .readdata
		.video_pixel_buffer_dma_0_avalon_control_slave_writedata        (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_writedata),  //                                                     .writedata
		.video_pixel_buffer_dma_0_avalon_control_slave_byteenable       (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_byteenable)  //                                                     .byteenable
	);

	oscill_nios_irq_mapper irq_mapper (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.sender_irq    (niosii_irq_irq)                      //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (audio_pll_reset_source_reset),   // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (pll_vga_outclk0_clk),                //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
