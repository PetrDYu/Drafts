// AUDIO_PLL.v

// Generated using ACDS version 16.0 211

`timescale 1 ps / 1 ps
module AUDIO_PLL (
		output wire  audio_pll_0_audio_clk_clk,      //    audio_pll_0_audio_clk.clk
		input  wire  audio_pll_0_ref_clk_clk,        //      audio_pll_0_ref_clk.clk
		input  wire  audio_pll_0_ref_reset_reset,    //    audio_pll_0_ref_reset.reset
		output wire  audio_pll_0_reset_source_reset  // audio_pll_0_reset_source.reset
	);

	AUDIO_PLL_audio_pll_0 audio_pll_0 (
		.ref_clk_clk        (audio_pll_0_ref_clk_clk),        //      ref_clk.clk
		.ref_reset_reset    (audio_pll_0_ref_reset_reset),    //    ref_reset.reset
		.audio_clk_clk      (audio_pll_0_audio_clk_clk),      //    audio_clk.clk
		.reset_source_reset (audio_pll_0_reset_source_reset)  // reset_source.reset
	);

endmodule
