// testVGAsystem.v

// Generated using ACDS version 16.0 211

`timescale 1 ps / 1 ps
module testVGAsystem (
		input  wire       clk_clk,                                         //                                       clk.clk
		input  wire       reset_reset_n,                                   //                                     reset.reset_n
		output wire       video_vga_controller_0_external_interface_CLK,   // video_vga_controller_0_external_interface.CLK
		output wire       video_vga_controller_0_external_interface_HS,    //                                          .HS
		output wire       video_vga_controller_0_external_interface_VS,    //                                          .VS
		output wire       video_vga_controller_0_external_interface_BLANK, //                                          .BLANK
		output wire       video_vga_controller_0_external_interface_SYNC,  //                                          .SYNC
		output wire [7:0] video_vga_controller_0_external_interface_R,     //                                          .R
		output wire [7:0] video_vga_controller_0_external_interface_G,     //                                          .G
		output wire [7:0] video_vga_controller_0_external_interface_B      //                                          .B
	);

	wire    pll_0_outclk0_clk;              // pll_0:outclk_0 -> [rst_controller:clk, video_vga_controller_0:clk]
	wire    rst_controller_reset_out_reset; // rst_controller:reset_out -> video_vga_controller_0:reset

	testVGAsystem_pll_0 pll_0 (
		.refclk   (clk_clk),           //  refclk.clk
		.rst      (~reset_reset_n),    //   reset.reset
		.outclk_0 (pll_0_outclk0_clk), // outclk0.clk
		.locked   ()                   // (terminated)
	);

	testVGAsystem_video_vga_controller_0 video_vga_controller_0 (
		.clk           (pll_0_outclk0_clk),                               //                clk.clk
		.reset         (rst_controller_reset_out_reset),                  //              reset.reset
		.data          (),                                                //    avalon_vga_sink.data
		.startofpacket (),                                                //                   .startofpacket
		.endofpacket   (),                                                //                   .endofpacket
		.valid         (),                                                //                   .valid
		.ready         (),                                                //                   .ready
		.VGA_CLK       (video_vga_controller_0_external_interface_CLK),   // external_interface.export
		.VGA_HS        (video_vga_controller_0_external_interface_HS),    //                   .export
		.VGA_VS        (video_vga_controller_0_external_interface_VS),    //                   .export
		.VGA_BLANK     (video_vga_controller_0_external_interface_BLANK), //                   .export
		.VGA_SYNC      (video_vga_controller_0_external_interface_SYNC),  //                   .export
		.VGA_R         (video_vga_controller_0_external_interface_R),     //                   .export
		.VGA_G         (video_vga_controller_0_external_interface_G),     //                   .export
		.VGA_B         (video_vga_controller_0_external_interface_B)      //                   .export
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (pll_0_outclk0_clk),              //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
